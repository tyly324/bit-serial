module decode